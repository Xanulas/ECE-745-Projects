package i2cmb_env_pkg;


import ncsu_pkg::*;
import i2c_pkg::*;
import wb_pkg::*;
import data_pkg::*;
`include "../../ncsu_pkg/ncsu_macros.svh"
`include "src/i2cmb_env_configuration.svh"
`include "src/i2cmb_generator.svh"
`include "src/i2cmb_scoreboard.svh"
`include "src/i2cmb_predictor.svh"
`include "src/i2cmb_coverage.svh"
`include "src/i2cmb_environment.svh"
`include "src/i2cmb_test.svh"

`include "src/test_i2cmb_consecutive_starts.svh"
`include "src/test_i2cmb_consecutive_stops.svh"
`include "src/test_i2cmb_reg_addr.svh"
`include "src/test_i2cmb_reg_vals.svh"   
`include "src/test_i2cmb_rw_ability.svh"        
`include "src/test_i2cmb_writes.svh"


endpackage