package wb_pkg;

import ncsu_pkg::*;
`include "../../ncsu_pkg/ncsu_macros.svh"
import data_pkg::*;
`include "src/wb_cfg.svh"
`include "src/wb_transaction.svh"
`include "src/wb_coverage.svh"
`include "src/wb_driver.svh"
`include "src/wb_monitor.svh"
`include "src/wb_agent.svh"

endpackage